
module Adder #(
    parameter BIT_WIDTH = 16)(
    input a,
    input b,
    output y);
endmodule
