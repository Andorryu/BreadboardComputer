
module top(
    
);
endmodule
